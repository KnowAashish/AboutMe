Hello World -GitHub
I want to push this file to GitHub.